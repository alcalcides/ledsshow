// by Alcides Augusto Bezerra Neto
// Turns led on and of
module ledsshow(led, pushButton);
	output led;
	input pushButton;
	
	assign led = pushButton;
	



endmodule